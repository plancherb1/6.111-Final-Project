// Switch Debounce Module
// use your system clock for the clock input
// to produce a synchronous, debounced output
// parameter: 27mhz clock: 270000, 25mhz clock: 250000 for .01 seconds
module debounce #(parameter DELAY=270000)
	        (input reset, clock, noisy,
	         output reg clean);

   reg [18:0] count;
   reg new;

   always @(posedge clock)
     if (reset)
       begin
	  count <= 0;
	  new <= noisy;
	  clean <= noisy;
       end
     else if (noisy != new)
       begin
	  new <= noisy;
	  count <= 0;
       end
     else if (count == DELAY)
       clean <= new;
     else
       count <= count+1;
      
endmodule