library verilog;
use verilog.vl_types.all;
entity main_fsm_tb is
end main_fsm_tb;
