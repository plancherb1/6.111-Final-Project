library verilog;
use verilog.vl_types.all;
entity median_5_tb is
end median_5_tb;
