library verilog;
use verilog.vl_types.all;
entity orientation_math_tb is
end orientation_math_tb;
