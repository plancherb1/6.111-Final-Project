library verilog;
use verilog.vl_types.all;
entity median_3_tb is
end median_3_tb;
