library verilog;
use verilog.vl_types.all;
entity find_min_5_vals_cascading_tb is
end find_min_5_vals_cascading_tb;
