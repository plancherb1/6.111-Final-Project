library verilog;
use verilog.vl_types.all;
entity calc_rsin_15_165_30_tb is
end calc_rsin_15_165_30_tb;
