//////////////////////////////////////////////////////////////////////////////////
// Company:        MIT 6.111 Final Project
// Engineer:       Brian Plancher
// 
// Module Name:    Ultrasound Location Calculator
// Project Name:   FPGA Phone Home
//
//////////////////////////////////////////////////////////////////////////////////

module ultrasound_location_calculator(
	input clock,
	input reset,
    input [11:0] ultrasound_signals,
    output reg done,
    output reg [11:0] rover_location,
	output reg [11:0] ultrasound_commands
	// output analyzer_clock, // for debug only
	// output [15:0] analyzer_data // for debug only
	);
	
	// TBD DO IT
	
endmodule	 